module bitboard (
);


    
endmodule